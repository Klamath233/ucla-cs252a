`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    19:40:18 04/15/2017 
// Design Name: 
// Module Name:    ppa 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module ppa(x, y, c_in, z, c_out);

parameter n;

input [15:0] x,
input [15:0] y,
input c_in,
output [15:0] z,
output c_out

wire
endmodule
